`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2025/05/21 23:27:34
// Design Name: 
// Module Name: SIM_uart_drive_TB
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module SIM_uart_drive_TB(

    );

reg    clk,rst    ;

initial begin
    rst = 1       ;
    #100          ;
    rst = 0       ;
    

end

always @() begin
    
end
endmodule
